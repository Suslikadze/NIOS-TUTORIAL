-- UART_NIOSII.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity UART_NIOSII is
	port (
		clk_clk       : in  std_logic := '0'; --    clk.clk
		reset_reset_n : in  std_logic := '0'; --  reset.reset_n
		serial_rxd    : in  std_logic := '0'; -- serial.rxd
		serial_txd    : out std_logic         --       .txd
	);
end entity UART_NIOSII;

architecture rtl of UART_NIOSII is
	component UART_NIOSII_HostPC is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(18 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(18 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component UART_NIOSII_HostPC;

	component UART_NIOSII_Memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component UART_NIOSII_Memory;

	component UART_NIOSII_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component UART_NIOSII_uart;

	component UART_NIOSII_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			HostPC_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			Memory_reset1_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			HostPC_data_master_address                : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			HostPC_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			HostPC_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			HostPC_data_master_read                   : in  std_logic                     := 'X';             -- read
			HostPC_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			HostPC_data_master_write                  : in  std_logic                     := 'X';             -- write
			HostPC_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			HostPC_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			HostPC_instruction_master_address         : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			HostPC_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			HostPC_instruction_master_read            : in  std_logic                     := 'X';             -- read
			HostPC_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			HostPC_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			HostPC_debug_mem_slave_write              : out std_logic;                                        -- write
			HostPC_debug_mem_slave_read               : out std_logic;                                        -- read
			HostPC_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HostPC_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			HostPC_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			HostPC_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			HostPC_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			Memory_s1_address                         : out std_logic_vector(14 downto 0);                    -- address
			Memory_s1_write                           : out std_logic;                                        -- write
			Memory_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Memory_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			Memory_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			Memory_s1_chipselect                      : out std_logic;                                        -- chipselect
			Memory_s1_clken                           : out std_logic;                                        -- clken
			uart_s1_address                           : out std_logic_vector(2 downto 0);                     -- address
			uart_s1_write                             : out std_logic;                                        -- write
			uart_s1_read                              : out std_logic;                                        -- read
			uart_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			uart_s1_begintransfer                     : out std_logic;                                        -- begintransfer
			uart_s1_chipselect                        : out std_logic                                         -- chipselect
		);
	end component UART_NIOSII_mm_interconnect_0;

	component UART_NIOSII_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component UART_NIOSII_irq_mapper;

	component uart_niosii_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component uart_niosii_rst_controller;

	component uart_niosii_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component uart_niosii_rst_controller_001;

	signal hostpc_data_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:HostPC_data_master_readdata -> HostPC:d_readdata
	signal hostpc_data_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:HostPC_data_master_waitrequest -> HostPC:d_waitrequest
	signal hostpc_data_master_debugaccess                       : std_logic;                     -- HostPC:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:HostPC_data_master_debugaccess
	signal hostpc_data_master_address                           : std_logic_vector(18 downto 0); -- HostPC:d_address -> mm_interconnect_0:HostPC_data_master_address
	signal hostpc_data_master_byteenable                        : std_logic_vector(3 downto 0);  -- HostPC:d_byteenable -> mm_interconnect_0:HostPC_data_master_byteenable
	signal hostpc_data_master_read                              : std_logic;                     -- HostPC:d_read -> mm_interconnect_0:HostPC_data_master_read
	signal hostpc_data_master_write                             : std_logic;                     -- HostPC:d_write -> mm_interconnect_0:HostPC_data_master_write
	signal hostpc_data_master_writedata                         : std_logic_vector(31 downto 0); -- HostPC:d_writedata -> mm_interconnect_0:HostPC_data_master_writedata
	signal hostpc_instruction_master_readdata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:HostPC_instruction_master_readdata -> HostPC:i_readdata
	signal hostpc_instruction_master_waitrequest                : std_logic;                     -- mm_interconnect_0:HostPC_instruction_master_waitrequest -> HostPC:i_waitrequest
	signal hostpc_instruction_master_address                    : std_logic_vector(18 downto 0); -- HostPC:i_address -> mm_interconnect_0:HostPC_instruction_master_address
	signal hostpc_instruction_master_read                       : std_logic;                     -- HostPC:i_read -> mm_interconnect_0:HostPC_instruction_master_read
	signal mm_interconnect_0_hostpc_debug_mem_slave_readdata    : std_logic_vector(31 downto 0); -- HostPC:debug_mem_slave_readdata -> mm_interconnect_0:HostPC_debug_mem_slave_readdata
	signal mm_interconnect_0_hostpc_debug_mem_slave_waitrequest : std_logic;                     -- HostPC:debug_mem_slave_waitrequest -> mm_interconnect_0:HostPC_debug_mem_slave_waitrequest
	signal mm_interconnect_0_hostpc_debug_mem_slave_debugaccess : std_logic;                     -- mm_interconnect_0:HostPC_debug_mem_slave_debugaccess -> HostPC:debug_mem_slave_debugaccess
	signal mm_interconnect_0_hostpc_debug_mem_slave_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:HostPC_debug_mem_slave_address -> HostPC:debug_mem_slave_address
	signal mm_interconnect_0_hostpc_debug_mem_slave_read        : std_logic;                     -- mm_interconnect_0:HostPC_debug_mem_slave_read -> HostPC:debug_mem_slave_read
	signal mm_interconnect_0_hostpc_debug_mem_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:HostPC_debug_mem_slave_byteenable -> HostPC:debug_mem_slave_byteenable
	signal mm_interconnect_0_hostpc_debug_mem_slave_write       : std_logic;                     -- mm_interconnect_0:HostPC_debug_mem_slave_write -> HostPC:debug_mem_slave_write
	signal mm_interconnect_0_hostpc_debug_mem_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:HostPC_debug_mem_slave_writedata -> HostPC:debug_mem_slave_writedata
	signal mm_interconnect_0_memory_s1_chipselect               : std_logic;                     -- mm_interconnect_0:Memory_s1_chipselect -> Memory:chipselect
	signal mm_interconnect_0_memory_s1_readdata                 : std_logic_vector(31 downto 0); -- Memory:readdata -> mm_interconnect_0:Memory_s1_readdata
	signal mm_interconnect_0_memory_s1_address                  : std_logic_vector(14 downto 0); -- mm_interconnect_0:Memory_s1_address -> Memory:address
	signal mm_interconnect_0_memory_s1_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Memory_s1_byteenable -> Memory:byteenable
	signal mm_interconnect_0_memory_s1_write                    : std_logic;                     -- mm_interconnect_0:Memory_s1_write -> Memory:write
	signal mm_interconnect_0_memory_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:Memory_s1_writedata -> Memory:writedata
	signal mm_interconnect_0_memory_s1_clken                    : std_logic;                     -- mm_interconnect_0:Memory_s1_clken -> Memory:clken
	signal mm_interconnect_0_uart_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	signal mm_interconnect_0_uart_s1_readdata                   : std_logic_vector(15 downto 0); -- uart:readdata -> mm_interconnect_0:uart_s1_readdata
	signal mm_interconnect_0_uart_s1_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_s1_address -> uart:address
	signal mm_interconnect_0_uart_s1_read                       : std_logic;                     -- mm_interconnect_0:uart_s1_read -> mm_interconnect_0_uart_s1_read:in
	signal mm_interconnect_0_uart_s1_begintransfer              : std_logic;                     -- mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	signal mm_interconnect_0_uart_s1_write                      : std_logic;                     -- mm_interconnect_0:uart_s1_write -> mm_interconnect_0_uart_s1_write:in
	signal mm_interconnect_0_uart_s1_writedata                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_s1_writedata -> uart:writedata
	signal irq_mapper_receiver0_irq                             : std_logic;                     -- uart:irq -> irq_mapper:receiver0_irq
	signal hostpc_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> HostPC:irq
	signal rst_controller_reset_out_reset                       : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:HostPC_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                   : std_logic;                     -- rst_controller:reset_req -> [HostPC:reset_req, rst_translator:reset_req_in]
	signal hostpc_debug_reset_request_reset                     : std_logic;                     -- HostPC:debug_reset_request -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                   : std_logic;                     -- rst_controller_001:reset_out -> [Memory:reset, mm_interconnect_0:Memory_reset1_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset_req               : std_logic;                     -- rst_controller_001:reset_req -> Memory:reset_req
	signal reset_reset_n_ports_inv                              : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_uart_s1_read_ports_inv             : std_logic;                     -- mm_interconnect_0_uart_s1_read:inv -> uart:read_n
	signal mm_interconnect_0_uart_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_uart_s1_write:inv -> uart:write_n
	signal rst_controller_reset_out_reset_ports_inv             : std_logic;                     -- rst_controller_reset_out_reset:inv -> [HostPC:reset_n, uart:reset_n]

begin

	hostpc : component UART_NIOSII_HostPC
		port map (
			clk                                 => clk_clk,                                              --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                           => hostpc_data_master_address,                           --               data_master.address
			d_byteenable                        => hostpc_data_master_byteenable,                        --                          .byteenable
			d_read                              => hostpc_data_master_read,                              --                          .read
			d_readdata                          => hostpc_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => hostpc_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => hostpc_data_master_write,                             --                          .write
			d_writedata                         => hostpc_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => hostpc_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => hostpc_instruction_master_address,                    --        instruction_master.address
			i_read                              => hostpc_instruction_master_read,                       --                          .read
			i_readdata                          => hostpc_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => hostpc_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => hostpc_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => hostpc_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_hostpc_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_hostpc_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_hostpc_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_hostpc_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_hostpc_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_hostpc_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_hostpc_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_hostpc_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                  -- custom_instruction_master.readra
		);

	memory : component UART_NIOSII_Memory
		port map (
			clk        => clk_clk,                                --   clk1.clk
			address    => mm_interconnect_0_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,     -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req, --       .reset_req
			freeze     => '0'                                     -- (terminated)
		);

	uart : component UART_NIOSII_uart
		port map (
			clk           => clk_clk,                                   --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_uart_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_s1_readdata,        --                    .readdata
			rxd           => serial_rxd,                                -- external_connection.export
			txd           => serial_txd,                                --                    .export
			irq           => irq_mapper_receiver0_irq                   --                 irq.irq
		);

	mm_interconnect_0 : component UART_NIOSII_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                              --                           clk_0_clk.clk
			HostPC_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                       --  HostPC_reset_reset_bridge_in_reset.reset
			Memory_reset1_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                   -- Memory_reset1_reset_bridge_in_reset.reset
			HostPC_data_master_address                => hostpc_data_master_address,                           --                  HostPC_data_master.address
			HostPC_data_master_waitrequest            => hostpc_data_master_waitrequest,                       --                                    .waitrequest
			HostPC_data_master_byteenable             => hostpc_data_master_byteenable,                        --                                    .byteenable
			HostPC_data_master_read                   => hostpc_data_master_read,                              --                                    .read
			HostPC_data_master_readdata               => hostpc_data_master_readdata,                          --                                    .readdata
			HostPC_data_master_write                  => hostpc_data_master_write,                             --                                    .write
			HostPC_data_master_writedata              => hostpc_data_master_writedata,                         --                                    .writedata
			HostPC_data_master_debugaccess            => hostpc_data_master_debugaccess,                       --                                    .debugaccess
			HostPC_instruction_master_address         => hostpc_instruction_master_address,                    --           HostPC_instruction_master.address
			HostPC_instruction_master_waitrequest     => hostpc_instruction_master_waitrequest,                --                                    .waitrequest
			HostPC_instruction_master_read            => hostpc_instruction_master_read,                       --                                    .read
			HostPC_instruction_master_readdata        => hostpc_instruction_master_readdata,                   --                                    .readdata
			HostPC_debug_mem_slave_address            => mm_interconnect_0_hostpc_debug_mem_slave_address,     --              HostPC_debug_mem_slave.address
			HostPC_debug_mem_slave_write              => mm_interconnect_0_hostpc_debug_mem_slave_write,       --                                    .write
			HostPC_debug_mem_slave_read               => mm_interconnect_0_hostpc_debug_mem_slave_read,        --                                    .read
			HostPC_debug_mem_slave_readdata           => mm_interconnect_0_hostpc_debug_mem_slave_readdata,    --                                    .readdata
			HostPC_debug_mem_slave_writedata          => mm_interconnect_0_hostpc_debug_mem_slave_writedata,   --                                    .writedata
			HostPC_debug_mem_slave_byteenable         => mm_interconnect_0_hostpc_debug_mem_slave_byteenable,  --                                    .byteenable
			HostPC_debug_mem_slave_waitrequest        => mm_interconnect_0_hostpc_debug_mem_slave_waitrequest, --                                    .waitrequest
			HostPC_debug_mem_slave_debugaccess        => mm_interconnect_0_hostpc_debug_mem_slave_debugaccess, --                                    .debugaccess
			Memory_s1_address                         => mm_interconnect_0_memory_s1_address,                  --                           Memory_s1.address
			Memory_s1_write                           => mm_interconnect_0_memory_s1_write,                    --                                    .write
			Memory_s1_readdata                        => mm_interconnect_0_memory_s1_readdata,                 --                                    .readdata
			Memory_s1_writedata                       => mm_interconnect_0_memory_s1_writedata,                --                                    .writedata
			Memory_s1_byteenable                      => mm_interconnect_0_memory_s1_byteenable,               --                                    .byteenable
			Memory_s1_chipselect                      => mm_interconnect_0_memory_s1_chipselect,               --                                    .chipselect
			Memory_s1_clken                           => mm_interconnect_0_memory_s1_clken,                    --                                    .clken
			uart_s1_address                           => mm_interconnect_0_uart_s1_address,                    --                             uart_s1.address
			uart_s1_write                             => mm_interconnect_0_uart_s1_write,                      --                                    .write
			uart_s1_read                              => mm_interconnect_0_uart_s1_read,                       --                                    .read
			uart_s1_readdata                          => mm_interconnect_0_uart_s1_readdata,                   --                                    .readdata
			uart_s1_writedata                         => mm_interconnect_0_uart_s1_writedata,                  --                                    .writedata
			uart_s1_begintransfer                     => mm_interconnect_0_uart_s1_begintransfer,              --                                    .begintransfer
			uart_s1_chipselect                        => mm_interconnect_0_uart_s1_chipselect                  --                                    .chipselect
		);

	irq_mapper : component UART_NIOSII_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => hostpc_irq_irq                  --    sender.irq
		);

	rst_controller : component uart_niosii_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => hostpc_debug_reset_request_reset,   -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component uart_niosii_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_uart_s1_read_ports_inv <= not mm_interconnect_0_uart_s1_read;

	mm_interconnect_0_uart_s1_write_ports_inv <= not mm_interconnect_0_uart_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of UART_NIOSII
