
module UART_NIOSII (
	clk_clk,
	reset_reset_n,
	serial_rxd,
	serial_txd);	

	input		clk_clk;
	input		reset_reset_n;
	input		serial_rxd;
	output		serial_txd;
endmodule
